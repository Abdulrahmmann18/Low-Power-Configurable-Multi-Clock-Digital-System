module RST_SYNC_tb ();

	////////////////////////////////// parameters declaration ///////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////////////
	parameter NUM_STAGES = 2;
	parameter CLK_PERIOD = 100;

	///////////////////////////////////// signals declaration ///////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////////////

	reg 				 CLK_tb;
	reg 				 RST_tb;
	wire 				 SYNC_RST_tb;

	//////////////////////////////////// clk generation block ///////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////////////
	initial begin
		CLK_tb = 1'b0;
		forever #(CLK_PERIOD/2) CLK_tb = ~CLK_tb;
	end

	////////////////////////////////////// DUT Instantiation ////////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////////////
	RST_SYNC DUT (
		.CLK(CLK_tb), .RST(RST_tb), .SYNC_RST(SYNC_RST_tb)
	);

	//////////////////////////////////////// test stimilus //////////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////////////
	
	initial begin
		RST_TASK();
		#1000
		$stop;

	end


	///////////////////////////////////// Tasks definations /////////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////////////
	task RST_TASK;
		begin
			RST_tb = 1'b0;
			#(2*CLK_PERIOD)
			RST_tb = 1'b1;
		end
	endtask






endmodule